module kmean

fn test_point_distance() {
    assert 1 == 1
}
